module Imm_Gen(
    input [31:0] inst,
    output reg [31:0] imm_out
);
    always @* begin
        case (inst[6:0])
            7'b0010011, 7'b0000011: // I-type
                imm_out = { {20{inst[31]}}, inst[31:20] };
            7'b0100011: // S-type
                imm_out = { {20{inst[31]}}, inst[31:25], inst[11:7] };
            7'b1100011: // B-type
                imm_out = { {19{inst[31]}}, inst[31], inst[7], inst[30:25], inst[11:8], 1'b0 };
            7'b1101111: // J-type (jal)
                imm_out = { {11{inst[31]}}, inst[31], inst[19:12], inst[20], inst[30:21], 1'b0 };
            7'b1100111: // jalr
                imm_out = { {20{inst[31]}}, inst[31:20] };
            default:
                imm_out = 0;
        endcase
    end
endmodule
